

library IEEE;
use IEEE.std_logic_1164.all;

package array2d is
  type array32_bit is array(31 downto 0, 31 downto 0) of std_logic;
end array2d;