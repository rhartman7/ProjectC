library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.all;

entity pc_plus_4 is
  port(
    a_input           :       in  std_logic_vector(31 downto 0);  
	s_reset :	in std_logic;                                
    o_output    :      out  std_logic_vector(31 downto 0));    
end pc_plus_4;

architecture structure of pc_plus_4 is

component ALU_32_bit
  	port(
		a_in  : in std_logic_vector(31 downto 0);
		b_in 	: in std_logic_vector(31 downto 0);
		op 	: in std_logic_vector(2 downto 0);
		add_sub : in std_logic;
		load_type : in std_logic;
		result_out : out std_logic_vector(31 downto 0);
		overflow : out std_logic;
		zero_out : out std_logic;
		c_out 	: out std_logic);
end component;



signal s_c_out, s_zero_out, s_overflow : std_logic;
signal s_output : std_logic_vector(31 downto 0);
begin
  adder: ALU_32_bit    -- Add branch target to PC value
    port map(
     		a_in  =>a_input,
		b_in   =>x"00000004",
		op 	  =>"101",
		add_sub  => '0',
		load_type   =>'0',
		result_out   =>s_output,
		overflow   =>s_overflow,
		zero_out   =>s_zero_out,
		c_out 	  =>s_c_out);

process (s_reset, s_output)
begin 
if (s_reset = '1' )then
o_output <= x"00000000";
else
o_output <= s_output;
end if;
end process;

end structure;