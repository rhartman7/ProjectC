library IEEE;
use IEEE.std_logic_1164.all;
use work.all;

-- This is an empty entity so we don't need to declare ports
entity tb_alu_mult_shift is
end tb_alu_mult_shift;

architecture behavior of tb_alu_mult_shift is

-- Declare the component we are going to instantiate
component alu_mult_shift
  	port(
		a_in  : in std_logic_vector(31 downto 0);
		b_in 	: in std_logic_vector(31 downto 0);
		op 	: in std_logic_vector(2 downto 0);
		add_sub : in std_logic;
		load_type : in std_logic;
		sel_shift_v: in std_logic;
		shift_amount : in std_logic_vector(4 downto 0);
		sel_srl_sll : in std_logic;
		sel_srl_sra : in std_logic;
		load_alu_shift_mult : in std_logic_vector(1 downto 0);
		result_out : out std_logic_vector(31 downto 0);
		overflow : out std_logic;
		zero_out : out std_logic;
		c_out 	: out std_logic);
end component;


-- Signals to connect to the struct_ones module
signal s_add_sub, s_load_type, s_sel_shift_v, s_sel_srl_sll, s_sel_srl_sra, s_overflow_out, s_zero_out, s_c_out : std_logic;
signal s_a_in, s_b_in, s_result_out : std_logic_vector(31 downto 0);
signal s_load_alu_shift_mult: std_logic_vector(1 downto 0);
signal s_op_in : std_logic_vector(2 downto 0);
signal s_shift_amount: std_logic_vector(4 downto 0);


begin

DUT: alu_mult_shift
  port map(
		a_in  => s_a_in,
		b_in 	 => s_b_in,
		op 	 => s_op_in,
		add_sub  => s_add_sub,
		load_type  => s_load_type,
		sel_shift_v => s_sel_shift_v,
		shift_amount => s_shift_amount,
		sel_srl_sll => s_sel_srl_sll,
		sel_srl_sra => s_sel_srl_sra,
		load_alu_shift_mult => s_load_alu_shift_mult,
		result_out => s_result_out,
		overflow  => s_overflow_out,
		zero_out  =>s_zero_out,
		c_out 	 => s_c_out);

 

  -- Remember, a process executes sequentially
  -- and then if not told to 'wait' loops back
  -- around
  tester : process


  begin


	--and
	s_a_in  <= x"FFFF0000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "000";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

	--or
	s_a_in  <= x"FFFF0000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "001";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

	--xor
	s_a_in  <= x"FFFF0000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "010";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;
	
--nand
	s_a_in  <= x"FFFF0000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "011";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

--nor
	s_a_in  <= x"FFFF0000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "100";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

--add
	s_a_in  <= x"FFFF0000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "101";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

--sub
	s_a_in  <= x"FFFF0000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "101";
	s_add_sub <= '1';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

--slt
	s_a_in  <= x"FFFF0000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

--slt
	s_a_in  <= x"00000000";
	s_b_in <= x"0000FFFF";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

--sltu	
	s_a_in  <= x"FFFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='1';
	s_load_alu_shift_mult <= "00";	
	wait for 100 ns;

--mult
	s_a_in  <= x"FFFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "10";	
	wait for 100 ns;

--sll
	s_a_in  <= x"FFFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "01";	
	s_sel_shift_v <= '0';
	s_shift_amount <= "00001";
	s_sel_srl_sll <= '1';
	s_sel_srl_sra <='0';
	wait for 100 ns;

--srl
	s_a_in  <= x"FFFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "01";	
	s_sel_shift_v <= '0';
	s_shift_amount <= "00001";
	s_sel_srl_sll <= '0';
	s_sel_srl_sra <='0';
	wait for 100 ns;

--sra shift in 1
	s_a_in  <= x"8FFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "01";	
	s_sel_shift_v <= '0';
	s_shift_amount <= "00001";
	s_sel_srl_sll <= '0';
	s_sel_srl_sra <='1';
	wait for 100 ns;

--sra shift in 0
	s_a_in  <= x"0FFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "01";	
	s_sel_shift_v <= '0';
	s_shift_amount <= "00001";
	s_sel_srl_sll <= '0';
	s_sel_srl_sra <='1';
	wait for 100 ns;

--srav
	s_a_in  <= x"8FFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "01";	
	s_sel_shift_v <= '1';
	s_shift_amount <= "00001";
	s_sel_srl_sll <= '0';
	s_sel_srl_sra <='1';
	wait for 100 ns;

--srlv
	s_a_in  <= x"FFFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "01";	
	s_sel_shift_v <= '1';
	s_shift_amount <= "00001";
	s_sel_srl_sll <= '0';
	s_sel_srl_sra <='0';
	wait for 100 ns;

--sllv
	s_a_in  <= x"FFFFFFFF";
	s_b_in <= x"00000000";
	s_op_in <= "110";
	s_add_sub <= '0';
	s_load_type <='0';
	s_load_alu_shift_mult <= "01";	
	s_sel_shift_v <= '1';
	s_shift_amount <= "00001";
	s_sel_srl_sll <= '1';
	s_sel_srl_sra <='0';
	wait for 100 ns;

  end process;
  
end behavior;
