library IEEE;
use IEEE.std_logic_1164.all;
use work.all;

entity eightto1mux_32 is
  port(
    input_0        :       in  std_logic_vector(31 downto 0);
    input_1       :        in  std_logic_vector(31 downto 0);
    input_2        :       in  std_logic_vector(31 downto 0);
    input_3        :       in  std_logic_vector(31 downto 0);
    input_4        :       in  std_logic_vector(31 downto 0);
    input_5        :       in  std_logic_vector(31 downto 0);
    input_6        :       in  std_logic_vector(31 downto 0);
    input_7        :       in  std_logic_vector(31 downto 0);
    sel3         :       in  std_logic_vector(2 downto 0);
    output       :       out std_logic_vector(31 downto 0));
    
end eightto1mux_32;


architecture structure of eightto1mux_32 is
  
begin
  
  with sel3 select
  
    output <= input_0    when "000",
              input_1    when "001",
              input_2    when "010",
              input_3    when "011",
              input_4    when "100",
              input_5    when "101",
              input_6    when "110",
              input_7    when "111",
          x"00000000"    when others;

end structure;
