library IEEE;
use IEEE.std_logic_1164.all;
use work.all;

entity alu_mult_shift is
  	port(
		a_in  : in std_logic_vector(31 downto 0);
		b_in 	: in std_logic_vector(31 downto 0);
		op 	: in std_logic_vector(2 downto 0);
		add_sub : in std_logic;
		load_type : in std_logic;
		sel_shift_v: in std_logic;
		shift_amount : in std_logic_vector(4 downto 0);
		sel_srl_sll : in std_logic;
		sel_srl_sra : in std_logic;
		load_alu_shift_mult : in std_logic_vector(1 downto 0);
		result_out : out std_logic_vector(31 downto 0);
		overflow : out std_logic;
		zero_out : out std_logic;
		c_out 	: out std_logic);
end alu_mult_shift;



architecture structure of alu_mult_shift is 

component Multiplier

  port (
    a_input       :       in  std_logic_vector(31 downto 0);
    b_input       :       in  std_logic_vector(31 downto 0);
    out_32        :       out std_logic_vector(31 downto 0));
end component;

component barrel_shifter_32
	
  	port(
		a_in  : in std_logic_vector(31 downto 0);
		sel : in std_logic_vector(4 downto 0);
		sel_srl_sll : in std_logic;
		sel_srl_sra : in std_logic;
		output 	: out std_logic_vector(31 downto 0));
end component;



component ALU_32_bit
  	port(
		a_in  : in std_logic_vector(31 downto 0);
		b_in 	: in std_logic_vector(31 downto 0);
		op 	: in std_logic_vector(2 downto 0);
		add_sub : in std_logic;
		load_type : in std_logic;
		result_out : out std_logic_vector(31 downto 0);
		overflow : out std_logic;
		zero_out : out std_logic;
		c_out 	: out std_logic);
end component;


component mux_21_n
	generic(N : integer := 32);
  	port(i_X  : in std_logic_vector(N-1 downto 0);
		i_Y: in std_logic_vector(N-1 downto 0);
		s_1 : in std_logic;
		o_Z : out std_logic_vector(N-1 downto 0));
end component;

component mux_4_1_32
	generic(N : integer := 32);
  	port(	i_00  : in std_logic_vector(N-1 downto 0);
		i_01  : in std_logic_vector(N-1 downto 0);
		i_10  : in std_logic_vector(N-1 downto 0);
		i_11  : in std_logic_vector(N-1 downto 0);
		sel : in std_logic_vector(1 downto 0);
		o_Z : out std_logic_vector(N-1 downto 0));
end component;

component mux_21_5_bit
	generic(N : integer := 5);
  	port(i_X  : in std_logic_vector(N-1 downto 0);
		i_Y: in std_logic_vector(N-1 downto 0);
		s_1 : in std_logic;
		o_Z : out std_logic_vector(N-1 downto 0));
end component;




signal s_alu_result_out, s_barrell_shifter_result_out, s_multiplier_out: std_logic_vector(31 downto 0);
signal s_shift_v_shift: std_logic_vector(4 downto 0);

begin

alu_32_i : ALU_32_bit
  port map(
		a_in  => a_in,
		b_in 	 => b_in,
		op 	 => op,
		add_sub  => add_sub,
		load_type  => load_type,
		result_out => s_alu_result_out,
		overflow  => overflow,
		zero_out  =>zero_out,
		c_out 	 => c_out);

shift_shift_v: mux_21_5_bit
	port MAP(i_X => shift_amount,
		i_Y => a_in(4 downto 0),
		s_1 =>sel_shift_v,
		o_Z  =>s_shift_v_shift);

barel_shifter : barrel_shifter_32
	port MAP(
		a_in => b_in,
		sel => s_shift_v_shift,
		sel_srl_sll => sel_srl_sll,
		sel_srl_sra => sel_srl_sra,
		output => s_barrell_shifter_result_out);

multi : Multiplier 
	port MAP (
   		 a_input  => a_in,
    		b_input => b_in,
    		out_32=> s_multiplier_out);

mux_4_1_32_i : mux_4_1_32
	port MAP (
		i_00 =>s_alu_result_out,
		i_01  => s_barrell_shifter_result_out,
		i_10 => s_multiplier_out,
		i_11  => x"00000000",
		sel => load_alu_shift_mult,
		o_Z => result_out);
end structure;


