library IEEE;
use IEEE.std_logic_1164.all;
use work.all;

entity bit_reversal is
  	port(	input  : in std_logic_vector( 31 downto 0);
		output : out std_logic_vector(31 downto 0));
end bit_reversal;

architecture structure of bit_reversal is 
 begin
output(0) <= input(31);
output(1) <= input(30);
output(2) <= input(29);
output(3) <= input(28);
output(4) <= input(27);
output(5) <= input(26);
output(6) <= input(25);
output(7) <= input(24);
output(8) <= input(23);
output(9) <= input(22);
output(10) <= input(21);
output(11) <= input(20);
output(12) <= input(19);
output(13) <= input(18);
output(14) <= input(17);
output(15) <= input(16);
output(16) <= input(15);
output(17) <= input(14);
output(18) <= input(13);
output(19) <= input(12);
output(20) <= input(11);
output(21) <= input(10);
output(22) <= input(9);
output(23) <= input(8);
output(24) <= input(7);
output(25) <= input(6);
output(26) <= input(5);
output(27) <= input(4);
output(28) <= input(3);
output(29) <= input(2);
output(30) <= input(1);
output(31) <= input(0);

end structure;